library verilog;
use verilog.vl_types.all;
entity state_automaton_vlg_vec_tst is
end state_automaton_vlg_vec_tst;
